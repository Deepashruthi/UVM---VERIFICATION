// Write pointer Handler
module wptr_handler #(parameter Ptr_Width = 3) 
  ( input logic wclk, wrst_n, w_en, 
   input logic [Ptr_Width:0] g_rptr_sync,
   output logic [Ptr_Width:0] b_wptr, g_wptr,
   output logic full);
  
  logic [Ptr_Width:0] b_wptr_next;
  logic [Ptr_Width:0] g_wptr_next;
  
  logic wfull;
  
  assign b_wptr_next = b_wptr +(w_en && !full);
  assign g_wptr_next = (b_wptr_next>>1)^b_wptr_next;
  
  always_ff @(posedge wclk or negedge wrst_n) begin
    if(!wrst_n) begin
      b_wptr <= 0;
      g_wptr <= 0;
      full <= 0;
    end
    else begin
      b_wptr <= b_wptr_next;
      g_wptr <= g_wptr_next;
      full <= wfull;
    end
  end
  
  assign wfull = (g_wptr_next == {~g_rptr_sync[Ptr_Width:Ptr_Width-1],g_rptr_sync[Ptr_Width-2:0]});
endmodule
