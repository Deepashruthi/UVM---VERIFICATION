// Interface
interface dff_if;
  logic clk;
  logic rst;
  logic d;
  logic q;
endinterface
